-- sukundy 1 misto
with second select
	cas3 <= "11111100" when "000000", -- 0
			"01100000" when "000001", -- 1
			"11011010" when "000010", -- 2
			"11110010" when "000011", -- 3
			"01100110" when "000100", -- 4
			"10110110" when "000101", -- 5
			"10111110" when "000110", -- 6
			"11100000" when "000111", -- 7
			"11111110" when "001000", -- 8
			"11110110" when "001001", -- 9
			"11111100" when "001010", -- 10
			"01100000" when "001011", -- 11
			"11011010" when "001100", -- 12
			"11110010" when "001101", -- 13
			"01100110" when "001110", -- 14
			"10110110" when "001111", -- 15
			"10111110" when "010000", -- 16
			"11100000" when "010001", -- 17
			"11111110" when "010010", -- 18
			"11110110" when "010011", -- 19
			"11111100" when "010100", -- 20
			"01100000" when "010101", -- 21
			"11011010" when "010110", -- 22
			"11110010" when "010111", -- 23
			"01100110" when "011000", -- 24
			"10110110" when "011001", -- 25
			"10111110" when "011010", -- 26
			"11100000" when "011011", -- 27
			"11111110" when "011100", -- 28
			"11110110" when "011101", -- 29
			"11111100" when "011110", -- 30
			"01100000" when "011111", -- 31
			"11011010" when "100000", -- 32
			"11110010" when "100001", -- 33
			"01100110" when "100010", -- 34
			"10110110" when "100011", -- 35
			"10111110" when "100100", -- 36
			"11100000" when "100101", -- 37
			"11111110" when "100110", -- 38
			"11110110" when "100111", -- 39
			"11111100" when "101000", -- 40
			"01100000" when "101001", -- 41
			"11011010" when "101010", -- 42
			"11110010" when "101011", -- 43
			"01100110" when "101100", -- 44
			"10110110" when "101101", -- 45
			"10111110" when "101110", -- 46
			"11100000" when "101111", -- 47
			"11111110" when "110000", -- 48
			"11110110" when "110001", -- 49
			"11111100" when "110010", -- 50
			"01100000" when "110011", -- 51
			"11011010" when "110100", -- 52
			"11110010" when "110101", -- 53
			"01100110" when "110110", -- 54
			"10110110" when "110111", -- 55
			"10111110" when "111000", -- 56
			"11100000" when "111001", -- 57
			"11111110" when "111010", -- 58
			"11110110" when "111011", -- 59
			"00000000" when others; 

-- sekundy 2 misto
with second select
	cas2 <= "11111100" when "000000", -- 0
			"11111100" when "000001", -- 1
			"11111100" when "000010", -- 2
			"11111100" when "000011", -- 3
			"11111100" when "000100", -- 4
			"11111100" when "000101", -- 5
			"11111100" when "000110", -- 6
			"11111100" when "000111", -- 7
			"11111100" when "001000", -- 8
			"11111100" when "001001", -- 9
			"01100000" when "001010", -- 10
			"01100000" when "001011", -- 11
			"01100000" when "001100", -- 12
			"01100000" when "001101", -- 13
			"01100000" when "001110", -- 14
			"01100000" when "001111", -- 15
			"01100000" when "010000", -- 16
			"01100000" when "010001", -- 17
			"01100000" when "010010", -- 18
			"01100000" when "010011", -- 19
			"11011010" when "010100", -- 20
			"11011010" when "010101", -- 21
			"11011010" when "010110", -- 22
			"11011010" when "010111", -- 23
			"11011010" when "011000", -- 24
			"11011010" when "011001", -- 25
			"11011010" when "011010", -- 26
			"11011010" when "011011", -- 27
			"11011010" when "011100", -- 28
			"11011010" when "011101", -- 29
			"11110010" when "011110", -- 30
			"11110010" when "011111", -- 31
			"11110010" when "100000", -- 32
			"11110010" when "100001", -- 33
			"11110010" when "100010", -- 34
			"11110010" when "100011", -- 35
			"11110010" when "100100", -- 36
			"11110010" when "100101", -- 37
			"11110010" when "100110", -- 38
			"11110010" when "100111", -- 39
			"01100110" when "101000", -- 40
			"01100110" when "101001", -- 41
			"01100110" when "101010", -- 42
			"01100110" when "101011", -- 43
			"01100110" when "101100", -- 44
			"01100110" when "101101", -- 45
			"01100110" when "101110", -- 46
			"01100110" when "101111", -- 47
			"01100110" when "110000", -- 48
			"01100110" when "110001", -- 49
			"10110110" when "110010", -- 50
			"10110110" when "110011", -- 51
			"10110110" when "110100", -- 52
			"10110110" when "110101", -- 53
			"10110110" when "110110", -- 54
			"10110110" when "110111", -- 55
			"10110110" when "111000", -- 56
			"10110110" when "111001", -- 57
			"10110110" when "111010", -- 58
			"10110110" when "111011", -- 59
			"00000000" when others; 


-- minuty 1 misto
with minut select
	cas1 <= "11111100" when "00000", -- 0
			"01100000" when "00001", -- 1
			"11011010" when "00010", -- 2
			"11110010" when "00011", -- 3
			"01100110" when "00100", -- 4
			"10110110" when "00101", -- 5
			"10111110" when "00110", -- 6
			"11100000" when "00111", -- 7
			"11111110" when "01000", -- 8
			"11110110" when "01001", -- 9
			"11111100" when "01010", -- 10
			"01100000" when "01011", -- 11
			"11011010" when "01100", -- 12
			"11110010" when "01101", -- 13
			"01100110" when "01110", -- 14
			"10110110" when "01111", -- 15
			"10111110" when "10000", -- 16
			"11100000" when "10001", -- 17
			"11111110" when "10010", -- 18
			"11110110" when "10011", -- 19
			"11111100" when "10100", -- 20
			"00000000" when others; 

-- minuty 2 misto
with minut select
	cas0 <= "11111100" when "00000", -- 0
			"11111100" when "00001", -- 1
			"11111100" when "00010", -- 2
			"11111100" when "00011", -- 3
			"11111100" when "00100", -- 4
			"11111100" when "00101", -- 5
			"11111100" when "00110", -- 6
			"11111100" when "00111", -- 7
			"11111100" when "01000", -- 8
			"11111100" when "01001", -- 9
			"01100000" when "01010", -- 10
			"01100000" when "01011", -- 11
			"01100000" when "01100", -- 12
			"01100000" when "01101", -- 13
			"01100000" when "01110", -- 14
			"01100000" when "01111", -- 15
			"01100000" when "10000", -- 16
			"01100000" when "10001", -- 17
			"01100000" when "10010", -- 18
			"01100000" when "10011", -- 19
			"11011010" when "10100", -- 20
			"00000000" when others; 

-- hoste body 1 misto
with hoste select
	b_host1 <= "11111100" when "000000", -- 0
			"01100000" when "000001", -- 1
			"11011010" when "000010", -- 2
			"11110010" when "000011", -- 3
			"01100110" when "000100", -- 4
			"10110110" when "000101", -- 5
			"10111110" when "000110", -- 6
			"11100000" when "000111", -- 7
			"11111110" when "001000", -- 8
			"11110110" when "001001", -- 9
			"11111100" when "001010", -- 10
			"01100000" when "001011", -- 11
			"11011010" when "001100", -- 12
			"11110010" when "001101", -- 13
			"01100110" when "001110", -- 14
			"10110110" when "001111", -- 15
			"10111110" when "010000", -- 16
			"11100000" when "010001", -- 17
			"11111110" when "010010", -- 18
			"11110110" when "010011", -- 19
			"11111100" when "010100", -- 20
			"01100000" when "010101", -- 21
			"11011010" when "010110", -- 22
			"11110010" when "010111", -- 23
			"01100110" when "011000", -- 24
			"10110110" when "011001", -- 25
			"10111110" when "011010", -- 26
			"11100000" when "011011", -- 27
			"11111110" when "011100", -- 28
			"11110110" when "011101", -- 29
			"11111100" when "011110", -- 30
			"01100000" when "011111", -- 31
			"11011010" when "100000", -- 32
			"11110010" when "100001", -- 33
			"01100110" when "100010", -- 34
			"10110110" when "100011", -- 35
			"10111110" when "100100", -- 36
			"11100000" when "100101", -- 37
			"11111110" when "100110", -- 38
			"11110110" when "100111", -- 39
			"11111100" when "101000", -- 40
			"01100000" when "101001", -- 41
			"11011010" when "101010", -- 42
			"11110010" when "101011", -- 43
			"01100110" when "101100", -- 44
			"10110110" when "101101", -- 45
			"10111110" when "101110", -- 46
			"11100000" when "101111", -- 47
			"11111110" when "110000", -- 48
			"11110110" when "110001", -- 49
			"11111100" when "110010", -- 50
			"01100000" when "110011", -- 51
			"11011010" when "110100", -- 52
			"11110010" when "110101", -- 53
			"01100110" when "110110", -- 54
			"10110110" when "110111", -- 55
			"10111110" when "111000", -- 56
			"11100000" when "111001", -- 57
			"11111110" when "111010", -- 58
			"11110110" when "111011", -- 59
			"00000000" when others; 